//
// Copyright 2021 Ziliang Guo
//
// Redistribution and use in source and binary forms, with or without modification,
// are permitted provided that the following conditions are met:
//
// 1. Redistributions of source code must retain the above copyright notice, this
// list of conditions and the following disclaimer.
// 2. Redistributions in binary form must reproduce the above copyright notice,
// this list of conditions and the following disclaimer in the documentation and/or
// other materials provided with the distribution.
// 3. Neither the name of the copyright holder nor the names of its contributors may
// be used to endorse or promote products derived from this software without specific
// prior written permission.
//
// THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS"
// AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE
// IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE
// ARE DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTORS BE
// LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR
// CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE
// GOODS OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION)
// HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT
// LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT
// OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
//

`timescale 1ns / 1ps

interface valid_intr();

  parameter int DATA_WIDTH = 32;

  logic [DATA_WIDTH-1:0] data;
  logic valid;

  modport master(
    output valid,
    output data
  );

  modport slave(
    input valid,
    input data
  );

endinterface

interface valid_burst_intr();

  parameter int DATA_WIDTH = 32;

  logic [DATA_WIDTH-1:0] data;
  logic valid;
  logic last;

  modport master(
    output valid,
    output last,
    output data
  );

  modport slave(
    input valid,
    output last,
    input data
  );

endinterface

interface decoupled_intr();

  parameter int DATA_WIDTH = 32;

  logic [DATA_WIDTH-1:0] data;
  logic valid;
  logic ready;

  modport master(
    output data,
    output valid,
    input ready
  );

  modport slave(
    input data,
    input valid,
    output ready
  );

endinterface

interface decoupled_burst_intr();

  parameter int DATA_WIDTH = 32;

  logic [DATA_WIDTH-1:0] data;
  logic valid;
  logic last;
  logic ready;

  modport master(
    output data,
    output valid,
    output last,
    input ready
  );

  modport slave(
    input data,
    input valid,
    input last,
    output ready
  );

endinterface
